-------------------------------------------------------------------
-- Arquivo   : comparador_85.vhd
-- Projeto   : Experiencia 2 - Um Fluxo de Dados Simples
-------------------------------------------------------------------
-- Descricao : comparador de magnitude de 4 bits 
--             similar ao CI 7485
--             baseado em descricao criada por Edson Gomi (11/2017)
-------------------------------------------------------------------
-- Revisoes  :
--     Data        Versao  Autor             Descricao
--     02/01/2021  1.0     Edson Midorikawa  criacao
--     07/01/2023  1.1     Edson Midorikawa  revisao
-------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity comparador_85 is
    port (
        i_A5   : in  std_logic;
        i_B5   : in  std_logic;
        i_A4   : in  std_logic;
        i_B4   : in  std_logic;
        i_A3   : in  std_logic;
        i_B3   : in  std_logic;
        i_A2   : in  std_logic;
        i_B2   : in  std_logic;
        i_A1   : in  std_logic;
        i_B1   : in  std_logic;
        i_A0   : in  std_logic;
        i_B0   : in  std_logic;
        i_AGTB : in  std_logic;
        i_ALTB : in  std_logic;
        i_AEQB : in  std_logic;
        o_AGTB : out std_logic;
        o_ALTB : out std_logic;
        o_AEQB : out std_logic
    );
end entity comparador_85;

architecture dataflow of comparador_85 is
    signal agtb : std_logic;
    signal aeqb : std_logic;
    signal altb : std_logic;
begin
  -- equacoes dos sinais: pagina 462, capitulo 6 do livro-texto
    -- Wakerly, J.F. Digital Design - Principles and Practice, 4th Edition
    -- veja tambem datasheet do CI SN7485 (Function Table) 
    agtb <= (i_A5 and not(i_B5)) or --Ver se A5 é maior que B5
            (not(i_A5 xor i_B5) and i_A4 and not(i_B4)) or --ver se A5 é igual a B5 e A4 é maior que B5
            (not(i_A5 xor i_B5) and not(i_A4 xor i_B4) and i_A3 and not(i_B3)) or --ver se A5 é igual a B5 e A4 é igual a B4 e A3 é maior que B3
            (not(i_A5 xor i_B5) and not(i_A4 xor i_B4) and not(i_A3 xor i_B3) and i_A2 and not(i_B2)) or --Repetir a lógica das linhas anteriores adicionando os sinais necessários
            (not(i_A5 xor i_B5) and not(i_A4 xor i_B4) and not(i_A3 xor i_B3) and not(i_A2 xor i_B2) and i_A1 and not(i_B1)) or
            (not(i_A5 xor i_B5) and not(i_A4 xor i_B4) and not(i_A3 xor i_B3) and not(i_A2 xor i_B2) and not(i_A1 xor i_B1) and i_A0 and not(i_B0));
    aeqb <= not((i_A5 xor i_B5) or (i_A4 xor i_B4) or (i_A3 xor i_B3) or (i_A2 xor i_B2) or (i_A1 xor i_B1) or (i_A0 xor i_B0));
    altb <= not(agtb or aeqb);
    -- saidas
    o_AGTB <= agtb or (aeqb and (not(i_AEQB) and not(i_ALTB)));
    o_ALTB <= altb or (aeqb and (not(i_AEQB) and not(i_AGTB)));
    o_AEQB <= aeqb and i_AEQB;
    
end architecture dataflow;

    
